
module InstructionMemory(Address, Instruction);
    input [31:0] Address;
    output reg [31:0] Instruction;
    
    always @(*)
        case (Address[31])
            1'b0:case (Address[9:2])
                8'd0:	Instruction<=32'b001000_00000_00100_00000_00000_000011;
                8'd1:	Instruction<=32'b001000_00100_00100_00000_00000_000001;
                8'd2:	Instruction<=32'b001000_00100_00100_00000_00000_000001;
                8'd3:	Instruction<=32'b001000_11101_11101_11111_11111_111100;
                8'd4:	Instruction<=32'b101011_11101_00100_00000_00000_000000;
                8'd5:	Instruction<=32'b100011_11101_00010_00000_00000_000000;
                8'd6:	Instruction<=32'b000100_00010_00100_00000_00000_000001;
                8'd7:	Instruction<=32'b000000_00010_00100_01000_00000_100000;
                8'd8:	Instruction<=32'b000000_01000_00010_01000_00000_100000;
                8'd9:	Instruction<=32'b000011_00000_00000_00000_00000_001010;
                8'd10:	Instruction<=32'b000000_00000_11111_00010_00000_100000;
                8'd11:	Instruction<=32'b100011_11101_01000_00000_00000_000000;
                8'd12:	Instruction<=32'b101011_11101_01000_11111_11111_111100;

                default: Instruction <= 32'h00000000;
            endcase
        1'b1:case (Address[9:2])
                8'd0:   Instruction<=32'b000010_00000_00000_00000_00000_000110;
                8'd1:   Instruction<=32'b000000_00000_00000_00000_00000_000000;
                8'd2:   Instruction<=32'b000010_00000_00000_00000_00000_000111;
                8'd3:   Instruction<=32'b000000_00000_00000_00000_00000_000000;
                8'd4:   Instruction<=32'b000010_00000_00000_00000_00000_001110;
                8'd5:   Instruction<=32'b000000_00000_00000_00000_00000_000000;
                8'd6:   Instruction<=32'b010000_10000_00000_00000_00000_011000;
                8'd7:   Instruction<=32'b100011_10000_11010_00000_00000_011000;
                8'd8:   Instruction<=32'b101011_11101_11010_00000_00000_000000;
                8'd9:   Instruction<=32'b101011_10000_00000_00000_00000_100000;
                8'd10:  Instruction<=32'b001000_11101_11101_00000_00000_000100;
                8'd11:  Instruction<=32'b001000_00000_00001_00000_00000_000001;
                8'd12:  Instruction<=32'b000000_00100_00001_00100_00000_100010;
                8'd13:  Instruction<=32'b010000_10000_00000_00000_00000_011000;
                8'd14:  Instruction<=32'b000010_00000_00000_00000_00000_001110;
                8'd15:  Instruction<=32'b000000_00000_00000_00000_00000_000000;                default: Instruction <= 32'h00000000;
            endcase
        endcase
endmodule
